module top_module (
    input in,
    output out);
wire w1;
    assign out = in;
endmodule
